class axi_lite_master_driver extends uvm_driver#(axi_lite_transaction);
	//Interface
	
